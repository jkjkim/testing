`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JT+31gRDptJqO+3i0+5tZMwsOwWlyUwFeZnqDXdlKuB+ImGI7mZjTTBNjB4kxw92EuPHhJc2lf4t
hQ47FEFvScB+yyp1h+qsWLZ1dyJIvwo0DrTtKk7MKx4jzY1adjPTareDB6i+YTUxM55elaku62c8
pzsadogzTWLTT7SqykRoCoRT8YS8Bsm53AoXmJ5WKtmS/GFq/wUnBgc0NIaheFD1me+isiXhQCyG
2lUyd17toO0wnjIxQjYJhk0Zc2GhrlfBHIsYB7slu0EG6qh+lSAyCQr/qPN5luKrdQVyq81IfMYD
0bM9p5twMF3wj5Ig5tpDtHeDMZHFjBNgZ+bX3A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YOsYqs0pDerC4EZodJW0nPUQx7gAivt4dT9rSP1+FVO+LdbFn77+RZkyD4WirOFhXeU9Rvk+YHTo
rie4n89Azq/WUiqJ6JwfReIeCEUGh5ZM/fnr47+Cnl1pnBUa4gx1f42Og3IiJW4+cvAwPH1xUngY
IiW0UZURcScx/CcVw4w=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
HrPt08LHFjdsa2aRHkx1lU2xlc3ZlVE2l+or2Bo8yFnBuwcOvTo0mghzG2dg+tfRo6g4qa1dnEmH
hVRxXMh1itzK2y2wZN7mq4X8xi29ZjnsrmiQAgQ2cPjzm3if8S3il0lOf9GFZu9IfKCw7fSaaHuM
6RZeXjDY/LpslP9NjWs=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hW3Ona5gsnRxbk32w/cEg1nRp8t3H2PJ4NKa9T30GXE3fWFEP1DRun0h9R89473yd4nDkCVTew5Y
ZgLjnCx9tQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2864)
`pragma protect data_block
sF9qiKXwsXXdVveDxN4/5SezwZet/FZC1OiAqYdoVjothronczGXKfIcnDs4vujNBxFXZQlCrjA2
BK676k/gkfMwiuaKKgeBF88pYjjW18Gf4EztnXHi4LOlklWi8B9AuRZ0YHsfEMgD9U3/Hy6j5HJU
CMfO637uww4IlvIfgxDoDnBJMmrjprkVLeoJaCuqtAH6eJMJhjJUNu9LRLtAw9rdw31irlB//I98
p3V7vPcxGlMvY4WWS2wZOMY32sRC1+OvbSWTqAn2aveTKimFVvKiC3TPnQxVCQYqmFs/75ErhLyz
PpkUvSUmqQsfvcZnXkiilimT8blNVM4QPGc8xR9O6ZhvW+QNlsORbkuKlGmCl2bxXrXH5OjMrjZD
bK7DoszmSjOjNEwkTnq+e2W56Re0HSq6EASiJosHDzROB/yHH+z9qJJ71D+jTNYl/V81Ue+FxKKP
S7qrb6XHOhVc76vFY7SxItInO/GdyVK026XRvhM7wOUNXfu9oa6EWj89eEOLn2MDT7k7WI4tEmCF
T+7MH7zfns5X3rLTkwE639b/IcNoNtqg2a1cfPHWGtGB2gyfFJ2QJLod7LGiJKwQUCtDcJWKtLfi
+0hKXDKo0WmAnHXU8LdwS2ypA8dE1b1c1dmJqx+NgWUsatE29MDmecBWKFcCTSuoWNX7t02sNBUL
HjLOtB/l6Rzc0/GQeYL+KcO1iDGKY4P3PltM4RZiXlwGZ5cISj8nTcw9E8KcxEqLppOxkkSKRIsc
8XW4UUGAWeC+ofCtBe6kKNoMAoxlIX1LFCZRikKxqiGZqLMwe53qJ0RhoFw7+e9Di9WV7XJgVKjf
5p5IZldW2bEsZFA6adta1bA23af79/bskzIiy0F+ozNAxHMfooZKE8KsD1Hh6ziRWg35mFCR30Sf
oy13pM/0HYOlUatcpwFa1uIllUTqsKTP+L3cKfnMtTFYy993Ox8Kp8/SWponWUkoaRjYPHN+22oR
+7VaTHdj8EdfdE8o9b87Y5xerU3j/0R1TMuOhkOat9+yAXNQgyCHqbBBuB4OC5Q6xewioe47Bz3h
0W7WBpDfhmux4K0em8owD9xl9/nvSzCKTh/oF8LxYQAlHwhIIlaIyT59nmbJtq1VUwBRhyAjNLhE
BODTCWUyn1spj9IcIcznHiTBgU+p2B2oUUM9fpA6jSCvUq9bIZ/3gmeG2ClkVmk+QzfLYj9JRaFU
b4TKwgW2FG3ZRwsXz12ribJvBc7VX2eRbFa3IoADxLyLYtqMtfAIwPX5S5UE5Oz5Y62HCrmNBCa9
DNtuCOPIHN0mn5/ica0fFjNblfUC2wSzEiPyihceV3Awb95xLpUG9Ofthyuog7qAAuNLhD99g+4J
5hzj2jBEL+maKX4Jbzg6h4Wyl7CPxXAIJkn9kn7TaaR0DaLQgAa2BXtbVpZrO0z2D0Y+qOavhQcV
sNFFvAxR0xPi5F1EwAhSCftCUv1KP811FVq/LUVQyUtPjbwfBb9KmMKCDL72YVOuGU1imeyL9xj7
HlFyACUIZGYUf5a3NsDIHlIocxAp2TjcUYC3MG/T8JnstqkPWwZtnkLcsuKq2PJiw+C3MvW6pZGu
8LXCDPq/nD1vxxYsV8709Z1c5xcMPPb07q9mC6JdtqkJrIqGuUMu244ZLs00l1lHYyu9vFhcao9D
GE0Zbg6TxizN1WKDC0Z+awvjutPGLiKWmxfdKhTeZrJZxEAMPkY96qoWiGs/Rn934ZuzJAbwpo5W
w27iCWKo2HKm5VvxI8RxXELTiXlo+qJfugS/4BKzLdWZxRwR+4u9ZOWymDUoqK9rR50Q6RmtT0DI
b7mty/aVKHxsEh4+JRgdJtblcFnRePihu82cBSpzGML4QgCrMw8f0Kx7PnRh+3PKMFaQsA1EnCzG
uzF4uHyKWl2XVwEPSyniGdNJK4RI2IfhbQh9eVQ7YNEHVC4alTcjSLrM9dM4rzyDU8TE488HiuR7
9SH03xLptyW/9NH2MXpkyusqIV2m+E9xEvCo02nBKiLd0909u4K8ZvrWYG2G7QZZE+p+5dvKrTzx
0Jngq3kdhSQNvp5AfKVkkxsOxKHcN6zjJTlWq/3ookGzqVHdlpbeN0kaeybIu1pUbchTM5WgNv5z
M0ZImpgQTFrFGJBUPR5htxsBFdxj3GP6oeZ8wifgAEn5AUkIpFG2ecWSziTDlcoZ4O/9Py7Icbnm
/9vdqsU9C2ociE4Oq7Bd3wwc7yds02G+DLYQ2HhGnRYiUdM2TrZJf/jeDeBAZvj836EF+7Dpcxv/
I6A34BttWmWhY+nI2D4F/mdDO/QejPUX6C1Cg9rIV+aUotGrHx2P5q2qA/HkqdPR1ceYR07npumo
NnhgDsFm48o835h+Kx3e2wctwnFuN1+uAI2oL2GQCoPBmTmNsb0WGIgE/mefcVovDbZAH7l2YD+p
zolqXyQfmJOtX5pwYaDIuEnVLSZpHf1+QKwfZHMae7AAPJp6XUwQBEaC8154TIrMcQH6619lIab0
/82ggDCCNJl2p1JaRiLNqdRbX1j/Qd7sVYcHbr2tMnY24oHTg9LofBxXK8pxB+yjKKK4Z/MIO1xt
kVe3c/+abRjJFS80Tg2kNwcsBZxQ7NYOQqgpn5bzcT8yZ7VN5VwHTt1JyLl4G+q0I6wkaaa7ppmZ
jNCIi+m6rv3lwtOkbDN9qzcIwn9SKnqlnfes6dQrWtnPO1MtbltBiLlAM1pWd4VP5HzVXoiQSn6k
4YZZshwNsIe6Sy7UFnOxuGOnC7oBzVWM1TQi7hnDeJpNJ3KsGAc4vsaZlH1y7IfpzUUxFg2AUaz8
wff90So8EIRh4CF08YhX/wNXaaoQO5YWcXTqCkt3Zm5cwRUSbDK9YMouVB4BV6G667c8RS8buLYi
GnkrKyPHttAMMlnajBbjXo151WRBFCZXV+6PwSh3iA0Mk2lJMlTKl3iZjh1zHBTcs+8KrBOEAruI
WiFEjj7xx+kAaVDtz2hQnqmi6IptN/D8Dm+FthwF0i2s8fUmpIFGEWrpXsFMRvdg7l9x5CvSGDYf
LwLUWWTYERRIIKZ+x1K8qgTjvSNRbcDW4dkLU9Yrs94Adph99viHaacAk/uvp1m0pWtIogvMY6R8
ok9bivVlEeX+KiCU2mzOSYHcoTlyTd+4h/zVd00Qm7LbIczOHE1CPCY4Ilk6gtEFlxy55AXz4jtS
0fJ/ZIszT79FLcNsT0r2vfrf17HbStbPX4QHNYMfkbstXF/i2Rm3wC+t8Obifbz4Ab48ZZMq3hTF
SUnclZl8f0/tSrz9TN2rRPu0UhEg3fHBgo0bTCdqkcCSDJvTWW/pS6J9rP8Q36vL07ESxqv7H3O7
JzvnMwRnkv/QKhlXl/YzPn1zlKadQ6yLUVZUEDMUv3dvyADaLGM1ExpGlGgPKf0PJNYDdz1OxYOM
Awiq1WF6hr6hFlmLadXvMzxWqNJiZXWYCZGMnOVvSBbEBScKZ0+N/2auiRtwUD6xbkGRkOxGKykz
XkT67D7zLhUiJxS+qQ3odcpT+gwlA+E+yzXnP+zwYC5qafPc0ZtReMjdFvH5DjkNEON6lKO8preT
+kSt8xPveV5QoXTJnZPEBX5q1iJQkQo36nzs6b0vRz57vO3h2lVyTSerHkyHzNf/MvHE7mLH8SI/
IgbZ92Q/BVi/A5uvEq04UbJQQDyOg1sThEafQ1wSKVflvZIskL/mdnS/PxEGPTOqRWcEkAudm4Y9
BRSRzQ8MWErT95F2VBIDF/fdPKYNseZa7J6xJdO+DQSmFPnBcZDKwT9FlrjpLmQ173p0Pw2pGxLB
3gYyXhwQ7PSlKocEbRU=
`pragma protect end_protected